if Instruction = "10111111" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10111111" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10111111" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10111111" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10111111" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10111111" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000000" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '1';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000001" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '1';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000010" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '1' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000101" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = '0' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = '1' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '1';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000100" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = '0' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000011" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='1';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000110" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '1';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10000111" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '1';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "11" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='0';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110001" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '1';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='0';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='0';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110000" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '0';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='0';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100000" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '1';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10100001" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '1';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '1';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '0';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110010" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '1';
                  MemWriteControl <= '0';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '0';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='0';

 elsif Instruction = "10110011" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '1';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10110011" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10110011" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10110011" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10110011" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '0';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10110011" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '0';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = '0' and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100010" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='1';
                  HighStackJump <= '0';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '0' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 1
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '1';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '1' and Q1 = '0' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '1' and Q1 = '1' and Q2 = '0' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '1';
                  InsRegControl <= '1';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '1' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '1';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '0' and Q1 = '1' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';

 elsif Instruction = "10100100" and Q0 = '0' and Q1 = '0' and Q2 = '1' and CarryFlag = 'X' and ABFlag = 'X' then
                  Count <= 0
                  CounterOutControl <= '0';
                  InsRegControl <= '0';
                  RegAControl <= '0';
                  RegBControl <= '0';
                  MainRegReadControl <= '0';
                  LowJumpRegLoad <= '0';
                  HighJumpRegLoad <= '0';
                  JumpEnable <= '0';
                  MainRegOutputControl <= '0';
                  MemOutEnable <= '0';
                  MemWriteControl <= '1';
                  Ram_LowControl <= '0';
                  Ram_HighControl <= '0';
                  Ram_Addr_Enable <='1';
                  StackCount <= '0';
                  StackOutControl <= '1';
                  DisplayControl <='0';
                  LowStackJump <='0';
                  HighStackJump <= '1';
                  StackCountDirection <='1';
else
                 Count <= 0
                 CounterOutControl <= '0';
                 InsRegControl <= '0';
                 RegAControl <= '0';
                 RegBControl <= '0';
                 MainRegReadControl <= '0';
                 LowJumpRegLoad <= '0';
                 HighJumpRegLoad <= '0';
                 JumpEnable <= '0';
                 MainRegOutputControl <= '1';
                 MemOutEnable <= '0';
                 MemWriteControl <= '1';
                 Ram_LowControl <= '0';
                 Ram_HighControl <= '0';
                 Ram_Addr_Enable <='1';
                 StackCount <= '0';
                 StackOutControl <= '1';
                 DisplayControl <='0';
                 LowStackJump <='0';
                 HighStackJump <= '0';
                 StackCountDirection <='1';
